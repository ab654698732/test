module m()
