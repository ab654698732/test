module m()
{}
